magic
tech sky130A
magscale 1 2
timestamp 1745686019
<< viali >>
rect 4997 9129 5031 9163
rect 5365 9061 5399 9095
rect 1409 8993 1443 9027
rect 1685 8925 1719 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 1593 8585 1627 8619
rect 1409 8449 1443 8483
rect 4445 8449 4479 8483
rect 4537 8449 4571 8483
rect 4261 8381 4295 8415
rect 4353 8313 4387 8347
rect 1409 7837 1443 7871
rect 5181 7837 5215 7871
rect 1593 7701 1627 7735
rect 5365 7701 5399 7735
rect 3341 7361 3375 7395
rect 3525 7361 3559 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 3433 7157 3467 7191
rect 4169 7157 4203 7191
rect 1409 6749 1443 6783
rect 5181 6749 5215 6783
rect 1593 6613 1627 6647
rect 5365 6613 5399 6647
rect 4721 6409 4755 6443
rect 3801 6273 3835 6307
rect 4537 6273 4571 6307
rect 3893 6205 3927 6239
rect 4169 6137 4203 6171
rect 3525 5865 3559 5899
rect 4077 5865 4111 5899
rect 1961 5729 1995 5763
rect 2237 5729 2271 5763
rect 3341 5729 3375 5763
rect 1869 5661 1903 5695
rect 3249 5661 3283 5695
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 3801 5593 3835 5627
rect 4261 5525 4295 5559
rect 1685 5185 1719 5219
rect 3157 5185 3191 5219
rect 5181 5185 5215 5219
rect 1409 5117 1443 5151
rect 3249 5117 3283 5151
rect 3525 5117 3559 5151
rect 5365 4981 5399 5015
rect 4353 4777 4387 4811
rect 3617 4709 3651 4743
rect 3341 4641 3375 4675
rect 3985 4641 4019 4675
rect 3249 4573 3283 4607
rect 4077 4573 4111 4607
rect 2513 4165 2547 4199
rect 1501 4097 1535 4131
rect 1777 4097 1811 4131
rect 1961 4097 1995 4131
rect 3801 4097 3835 4131
rect 3985 4097 4019 4131
rect 4261 4097 4295 4131
rect 5181 4097 5215 4131
rect 2053 4029 2087 4063
rect 4169 4029 4203 4063
rect 2513 3961 2547 3995
rect 4077 3961 4111 3995
rect 1685 3893 1719 3927
rect 5365 3893 5399 3927
rect 1593 3689 1627 3723
rect 1409 3485 1443 3519
rect 4445 3145 4479 3179
rect 5089 3145 5123 3179
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 4629 3009 4663 3043
rect 4721 3009 4755 3043
rect 4905 3009 4939 3043
rect 5273 3009 5307 3043
rect 5365 3009 5399 3043
rect 5089 2941 5123 2975
rect 4261 2873 4295 2907
rect 4813 2873 4847 2907
rect 1961 2601 1995 2635
rect 1685 2533 1719 2567
rect 1777 2397 1811 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 1501 2329 1535 2363
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 842 8984 848 9036
rect 900 9024 906 9036
rect 1397 9027 1455 9033
rect 1397 9024 1409 9027
rect 900 8996 1409 9024
rect 900 8984 906 8996
rect 1397 8993 1409 8996
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 4062 8956 4068 8968
rect 1719 8928 4068 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 3510 8848 3516 8900
rect 3568 8888 3574 8900
rect 5184 8888 5212 8919
rect 3568 8860 5212 8888
rect 3568 8848 3574 8860
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1627 8588 4568 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 4540 8492 4568 8588
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4062 8480 4068 8492
rect 3844 8452 4068 8480
rect 3844 8440 3850 8452
rect 4062 8440 4068 8452
rect 4120 8480 4126 8492
rect 4433 8483 4491 8489
rect 4433 8480 4445 8483
rect 4120 8452 4445 8480
rect 4120 8440 4126 8452
rect 4433 8449 4445 8452
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4522 8440 4528 8492
rect 4580 8440 4586 8492
rect 4246 8372 4252 8424
rect 4304 8372 4310 8424
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 4614 8344 4620 8356
rect 4387 8316 4620 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4488 7840 5181 7868
rect 4488 7828 4494 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 3878 7732 3884 7744
rect 1627 7704 3884 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 4246 7460 4252 7472
rect 3528 7432 4252 7460
rect 3528 7401 3556 7432
rect 4246 7420 4252 7432
rect 4304 7460 4310 7472
rect 5074 7460 5080 7472
rect 4304 7432 5080 7460
rect 4304 7420 4310 7432
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 3344 7256 3372 7355
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 4120 7364 4169 7392
rect 4120 7352 4126 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 4356 7324 4384 7355
rect 3752 7296 4384 7324
rect 3752 7284 3758 7296
rect 4706 7256 4712 7268
rect 3344 7228 4712 7256
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 3970 7188 3976 7200
rect 3467 7160 3976 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4154 7148 4160 7200
rect 4212 7148 4218 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 4212 6752 5181 6780
rect 4212 6740 4218 6752
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 3142 6644 3148 6656
rect 1627 6616 3148 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 4798 6440 4804 6452
rect 4755 6412 4804 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 4062 6304 4068 6316
rect 3835 6276 4068 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4798 6236 4804 6248
rect 3927 6208 4804 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4157 6171 4215 6177
rect 4157 6137 4169 6171
rect 4203 6168 4215 6171
rect 5166 6168 5172 6180
rect 4203 6140 5172 6168
rect 4203 6137 4215 6140
rect 4157 6131 4215 6137
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4706 6100 4712 6112
rect 4396 6072 4712 6100
rect 4396 6060 4402 6072
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 3510 5856 3516 5908
rect 3568 5856 3574 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3786 5896 3792 5908
rect 3660 5868 3792 5896
rect 3660 5856 3666 5868
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3844 5868 4077 5896
rect 3844 5856 3850 5868
rect 4065 5865 4077 5868
rect 4111 5896 4123 5899
rect 4890 5896 4896 5908
rect 4111 5868 4896 5896
rect 4111 5865 4123 5868
rect 4065 5859 4123 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 4614 5828 4620 5840
rect 3344 5800 4620 5828
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 1854 5652 1860 5704
rect 1912 5652 1918 5704
rect 1964 5692 1992 5723
rect 2222 5720 2228 5772
rect 2280 5720 2286 5772
rect 3344 5769 3372 5800
rect 4614 5788 4620 5800
rect 4672 5788 4678 5840
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 3050 5692 3056 5704
rect 1964 5664 3056 5692
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3602 5692 3608 5704
rect 3283 5664 3608 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3936 5664 3985 5692
rect 3936 5652 3942 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4246 5692 4252 5704
rect 4111 5664 4252 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 3142 5584 3148 5636
rect 3200 5624 3206 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 3200 5596 3801 5624
rect 3200 5584 3206 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 3234 5516 3240 5568
rect 3292 5556 3298 5568
rect 3988 5556 4016 5655
rect 4246 5652 4252 5664
rect 4304 5692 4310 5704
rect 4522 5692 4528 5704
rect 4304 5664 4528 5692
rect 4304 5652 4310 5664
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 3292 5528 4016 5556
rect 4249 5559 4307 5565
rect 3292 5516 3298 5528
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4338 5556 4344 5568
rect 4295 5528 4344 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4338 5516 4344 5528
rect 4396 5556 4402 5568
rect 4982 5556 4988 5568
rect 4396 5528 4988 5556
rect 4396 5516 4402 5528
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 3878 5284 3884 5296
rect 1688 5256 3884 5284
rect 1688 5225 1716 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 3142 5176 3148 5228
rect 3200 5176 3206 5228
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4396 5188 5181 5216
rect 4396 5176 4402 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 842 5108 848 5160
rect 900 5148 906 5160
rect 1397 5151 1455 5157
rect 1397 5148 1409 5151
rect 900 5120 1409 5148
rect 900 5108 906 5120
rect 1397 5117 1409 5120
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 4154 5148 4160 5160
rect 3559 5120 4160 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3252 5080 3280 5111
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4430 5080 4436 5092
rect 3252 5052 4436 5080
rect 4430 5040 4436 5052
rect 4488 5040 4494 5092
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 4338 4768 4344 4820
rect 4396 4768 4402 4820
rect 3605 4743 3663 4749
rect 3605 4709 3617 4743
rect 3651 4740 3663 4743
rect 4522 4740 4528 4752
rect 3651 4712 4528 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3234 4564 3240 4616
rect 3292 4564 3298 4616
rect 3344 4536 3372 4635
rect 3970 4632 3976 4684
rect 4028 4632 4034 4684
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3936 4576 4077 4604
rect 3936 4564 3942 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4706 4536 4712 4548
rect 3344 4508 4712 4536
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 2501 4199 2559 4205
rect 2501 4165 2513 4199
rect 2547 4196 2559 4199
rect 4154 4196 4160 4208
rect 2547 4168 4160 4196
rect 2547 4165 2559 4168
rect 2501 4159 2559 4165
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1535 4100 1777 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4128 2007 4131
rect 1995 4100 3004 4128
rect 1995 4097 2007 4100
rect 1949 4091 2007 4097
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 1964 4060 1992 4091
rect 1728 4032 1992 4060
rect 1728 4020 1734 4032
rect 2038 4020 2044 4072
rect 2096 4020 2102 4072
rect 2976 4060 3004 4100
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 3108 4100 3801 4128
rect 3108 4088 3114 4100
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4080 4100 4261 4128
rect 4080 4060 4108 4100
rect 4249 4097 4261 4100
rect 4295 4128 4307 4131
rect 4338 4128 4344 4140
rect 4295 4100 4344 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4338 4088 4344 4100
rect 4396 4128 4402 4140
rect 5074 4128 5080 4140
rect 4396 4100 5080 4128
rect 4396 4088 4402 4100
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 2976 4032 4108 4060
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4982 4060 4988 4072
rect 4212 4032 4988 4060
rect 4212 4020 4218 4032
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 1912 3964 2513 3992
rect 1912 3952 1918 3964
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 3712 3964 4016 3992
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 3712 3924 3740 3964
rect 1719 3896 3740 3924
rect 3988 3924 4016 3964
rect 4062 3952 4068 4004
rect 4120 3952 4126 4004
rect 5074 3924 5080 3936
rect 3988 3896 5080 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 4062 3720 4068 3732
rect 1627 3692 4068 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 842 3476 848 3528
rect 900 3516 906 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 900 3488 1409 3516
rect 900 3476 906 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 4430 3136 4436 3188
rect 4488 3136 4494 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 4580 3148 4752 3176
rect 4580 3136 4586 3148
rect 4724 3108 4752 3148
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 4856 3148 5089 3176
rect 4856 3136 4862 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 4264 3080 4660 3108
rect 4724 3080 4936 3108
rect 4264 3052 4292 3080
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4246 3040 4252 3052
rect 4203 3012 4252 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 4632 3049 4660 3080
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 4798 3040 4804 3052
rect 4755 3012 4804 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 4908 3049 4936 3080
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 4908 2972 4936 3003
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5040 3012 5273 3040
rect 5040 3000 5046 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 3292 2944 4844 2972
rect 4908 2944 5089 2972
rect 3292 2932 3298 2944
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2904 4307 2907
rect 4614 2904 4620 2916
rect 4295 2876 4620 2904
rect 4295 2873 4307 2876
rect 4249 2867 4307 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 4816 2913 4844 2944
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 4801 2907 4859 2913
rect 4801 2873 4813 2907
rect 4847 2873 4859 2907
rect 4801 2867 4859 2873
rect 3970 2796 3976 2848
rect 4028 2836 4034 2848
rect 5368 2836 5396 3003
rect 4028 2808 5396 2836
rect 4028 2796 4034 2808
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1854 2592 1860 2644
rect 1912 2632 1918 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 1912 2604 1961 2632
rect 1912 2592 1918 2604
rect 1949 2601 1961 2604
rect 1995 2601 2007 2635
rect 1949 2595 2007 2601
rect 1670 2524 1676 2576
rect 1728 2524 1734 2576
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 992 2400 1777 2428
rect 992 2388 998 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 1486 2320 1492 2372
rect 1544 2320 1550 2372
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 848 8984 900 9036
rect 4068 8916 4120 8968
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 3516 8848 3568 8900
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 3792 8440 3844 8492
rect 4068 8440 4120 8492
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 4620 8304 4672 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 848 7828 900 7880
rect 4436 7828 4488 7880
rect 3884 7692 3936 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 4252 7420 4304 7472
rect 5080 7420 5132 7472
rect 4068 7352 4120 7404
rect 3700 7284 3752 7336
rect 4712 7216 4764 7268
rect 3976 7148 4028 7200
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 848 6740 900 6792
rect 4160 6740 4212 6792
rect 3148 6604 3200 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 4804 6400 4856 6452
rect 4068 6264 4120 6316
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4804 6196 4856 6248
rect 5172 6128 5224 6180
rect 4344 6060 4396 6112
rect 4712 6060 4764 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 3608 5856 3660 5908
rect 3792 5856 3844 5908
rect 4896 5856 4948 5908
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 4620 5788 4672 5840
rect 3056 5652 3108 5704
rect 3608 5652 3660 5704
rect 3884 5652 3936 5704
rect 3148 5584 3200 5636
rect 3240 5516 3292 5568
rect 4252 5652 4304 5704
rect 4528 5652 4580 5704
rect 4344 5516 4396 5568
rect 4988 5516 5040 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 3884 5244 3936 5296
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 4344 5176 4396 5228
rect 848 5108 900 5160
rect 4160 5108 4212 5160
rect 4436 5040 4488 5092
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 4528 4700 4580 4752
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 3976 4675 4028 4684
rect 3976 4641 3985 4675
rect 3985 4641 4019 4675
rect 4019 4641 4028 4675
rect 3976 4632 4028 4641
rect 3884 4564 3936 4616
rect 4712 4496 4764 4548
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 4160 4156 4212 4208
rect 1676 4020 1728 4072
rect 2044 4063 2096 4072
rect 2044 4029 2053 4063
rect 2053 4029 2087 4063
rect 2087 4029 2096 4063
rect 2044 4020 2096 4029
rect 3056 4088 3108 4140
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4344 4088 4396 4140
rect 5080 4088 5132 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 4988 4020 5040 4072
rect 1860 3952 1912 4004
rect 4068 3995 4120 4004
rect 4068 3961 4077 3995
rect 4077 3961 4111 3995
rect 4111 3961 4120 3995
rect 4068 3952 4120 3961
rect 5080 3884 5132 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 4068 3680 4120 3732
rect 848 3476 900 3528
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 4436 3179 4488 3188
rect 4436 3145 4445 3179
rect 4445 3145 4479 3179
rect 4479 3145 4488 3179
rect 4436 3136 4488 3145
rect 4528 3136 4580 3188
rect 4804 3136 4856 3188
rect 4252 3000 4304 3052
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 4804 3000 4856 3052
rect 3240 2932 3292 2984
rect 4988 3000 5040 3052
rect 4620 2864 4672 2916
rect 3976 2796 4028 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 1860 2592 1912 2644
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 940 2388 992 2440
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 1492 2363 1544 2372
rect 1492 2329 1501 2363
rect 1501 2329 1535 2363
rect 1535 2329 1544 2363
rect 1492 2320 1544 2329
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 848 9036 900 9042
rect 848 8978 900 8984
rect 860 8945 888 8978
rect 846 8936 902 8945
rect 846 8871 902 8880
rect 1412 8498 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 5354 9007 5410 9016
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 848 7880 900 7886
rect 846 7848 848 7857
rect 900 7848 902 7857
rect 846 7783 902 7792
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 846 6488 902 6497
rect 2610 6491 2918 6500
rect 846 6423 902 6432
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 1860 5704 1912 5710
rect 2240 5681 2268 5714
rect 3056 5704 3108 5710
rect 1860 5646 1912 5652
rect 2226 5672 2282 5681
rect 848 5160 900 5166
rect 846 5128 848 5137
rect 900 5128 902 5137
rect 846 5063 902 5072
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 848 3528 900 3534
rect 846 3496 848 3505
rect 900 3496 902 3505
rect 846 3431 902 3440
rect 1688 2582 1716 4014
rect 1872 4010 1900 5646
rect 3056 5646 3108 5652
rect 2226 5607 2282 5616
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 3068 4146 3096 5646
rect 3160 5642 3188 6598
rect 3528 5914 3556 8842
rect 4080 8498 4108 8910
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3620 5710 3648 5850
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3160 5234 3188 5578
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3712 5522 3740 7278
rect 3804 5914 3832 8434
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3896 5710 3924 7686
rect 4264 7478 4292 8366
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3252 4622 3280 5510
rect 3712 5494 3924 5522
rect 3896 5302 3924 5494
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3896 4622 3924 5238
rect 3988 4690 4016 7142
rect 4080 6322 4108 7346
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 7041 4200 7142
rect 4158 7032 4214 7041
rect 4158 6967 4214 6976
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3884 4616 3936 4622
rect 3936 4564 4016 4570
rect 3884 4558 4016 4564
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2044 4072 2096 4078
rect 2042 4040 2044 4049
rect 2096 4040 2098 4049
rect 1860 4004 1912 4010
rect 2042 3975 2098 3984
rect 1860 3946 1912 3952
rect 1872 2650 1900 3946
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3252 2990 3280 4558
rect 3896 4542 4016 4558
rect 3988 4146 4016 4542
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3988 2854 4016 4082
rect 4080 4010 4108 6258
rect 4172 5166 4200 6734
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4172 4078 4200 4150
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4080 3738 4108 3946
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4264 3058 4292 5646
rect 4356 5574 4384 6054
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4448 5250 4476 7822
rect 4540 6322 4568 8434
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4540 5710 4568 6258
rect 4632 5930 4660 8298
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4724 6118 4752 7210
rect 4816 6458 4844 8910
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4632 5902 4752 5930
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4344 5228 4396 5234
rect 4448 5222 4568 5250
rect 4344 5170 4396 5176
rect 4356 4826 4384 5170
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4356 3074 4384 4082
rect 4448 3194 4476 5034
rect 4540 4758 4568 5222
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4540 3074 4568 3130
rect 4356 3058 4568 3074
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4344 3052 4568 3058
rect 4396 3046 4568 3052
rect 4344 2994 4396 3000
rect 4632 2922 4660 5782
rect 4724 4554 4752 5902
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4816 3194 4844 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4908 3074 4936 5850
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 4078 5028 5510
rect 5092 4146 5120 7414
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6361 5396 6598
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5184 4146 5212 6122
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 4816 3058 4936 3074
rect 5000 3058 5028 4014
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4804 3052 4936 3058
rect 4856 3046 4936 3052
rect 4988 3052 5040 3058
rect 4804 2994 4856 3000
rect 4988 2994 5040 3000
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 4618 2544 4674 2553
rect 4618 2479 4674 2488
rect 4632 2446 4660 2479
rect 5092 2446 5120 3878
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 952 2281 980 2382
rect 1492 2372 1544 2378
rect 1492 2314 1544 2320
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 938 2272 994 2281
rect 938 2207 994 2216
rect 1504 921 1532 2314
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1490 912 1546 921
rect 1490 847 1546 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 846 8880 902 8936
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 846 7828 848 7848
rect 848 7828 900 7848
rect 900 7828 902 7848
rect 846 7792 902 7828
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 846 6432 902 6488
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 846 5108 848 5128
rect 848 5108 900 5128
rect 900 5108 902 5128
rect 846 5072 902 5108
rect 846 3476 848 3496
rect 848 3476 900 3496
rect 900 3476 902 3496
rect 846 3440 902 3476
rect 2226 5616 2282 5672
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 4158 6976 4214 7032
rect 2042 4020 2044 4040
rect 2044 4020 2096 4040
rect 2096 4020 2098 4040
rect 2042 3984 2098 4020
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 4618 2488 4674 2544
rect 5354 3576 5410 3632
rect 938 2216 994 2272
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1490 856 1546 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7850 907 7853
rect 798 7848 907 7850
rect 798 7792 846 7848
rect 902 7792 907 7848
rect 798 7787 907 7792
rect 798 7744 858 7787
rect 0 7654 858 7744
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 0 7624 800 7654
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 4153 7036 4219 7037
rect 4102 7034 4108 7036
rect 4062 6974 4108 7034
rect 4172 7032 4219 7036
rect 4214 6976 4219 7032
rect 4102 6972 4108 6974
rect 4172 6972 4219 6976
rect 4153 6971 4219 6972
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2221 5674 2287 5677
rect 4470 5674 4476 5676
rect 2221 5672 4476 5674
rect 2221 5616 2226 5672
rect 2282 5616 4476 5672
rect 2221 5614 4476 5616
rect 2221 5611 2287 5614
rect 4470 5612 4476 5614
rect 4540 5612 4546 5676
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 2037 4042 2103 4045
rect 4102 4042 4108 4044
rect 2037 4040 4108 4042
rect 2037 3984 2042 4040
rect 2098 3984 4108 4040
rect 2037 3982 4108 3984
rect 2037 3979 2103 3982
rect 4102 3980 4108 3982
rect 4172 3980 4178 4044
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 0 3634 800 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 0 3544 858 3634
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 798 3501 858 3544
rect 798 3496 907 3501
rect 798 3440 846 3496
rect 902 3440 907 3496
rect 798 3438 907 3440
rect 841 3435 907 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 4470 2484 4476 2548
rect 4540 2546 4546 2548
rect 4613 2546 4679 2549
rect 4540 2544 4679 2546
rect 4540 2488 4618 2544
rect 4674 2488 4679 2544
rect 4540 2486 4679 2488
rect 4540 2484 4546 2486
rect 4613 2483 4679 2486
rect 0 2274 800 2304
rect 933 2274 999 2277
rect 0 2272 999 2274
rect 0 2216 938 2272
rect 994 2216 999 2272
rect 0 2214 999 2216
rect 0 2184 800 2214
rect 933 2211 999 2214
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1485 914 1551 917
rect 0 912 1551 914
rect 0 856 1490 912
rect 1546 856 1551 912
rect 0 854 1551 856
rect 0 824 800 854
rect 1485 851 1551 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 4108 7032 4172 7036
rect 4108 6976 4158 7032
rect 4158 6976 4172 7032
rect 4108 6972 4172 6976
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 4476 5612 4540 5676
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 4108 3980 4172 4044
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 4476 2484 4540 2548
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 4107 7036 4173 7037
rect 4107 6972 4108 7036
rect 4172 6972 4173 7036
rect 4107 6971 4173 6972
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 4110 4045 4170 6971
rect 4475 5676 4541 5677
rect 4475 5612 4476 5676
rect 4540 5612 4541 5676
rect 4475 5611 4541 5612
rect 4107 4044 4173 4045
rect 4107 3980 4108 4044
rect 4172 3980 4173 4044
rect 4107 3979 4173 3980
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 4478 2549 4538 5611
rect 4475 2548 4541 2549
rect 4475 2484 4476 2548
rect 4540 2484 4541 2548
rect 4475 2483 4541 2484
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__nand2_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _12_
timestamp 1704896540
transform 1 0 3036 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _16_
timestamp 1704896540
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _17_
timestamp 1704896540
transform 1 0 3864 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _18_
timestamp 1704896540
transform -1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _20_
timestamp 1704896540
transform 1 0 3772 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _21_
timestamp 1704896540
transform 1 0 1656 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2668 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1704896540
transform -1 0 4784 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2024 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_47
timestamp 1704896540
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 1704896540
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18
timestamp 1704896540
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 1704896540
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_17
timestamp 1704896540
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_36
timestamp 1704896540
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_37
timestamp 1704896540
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_13
timestamp 1704896540
transform 1 0 2300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_19
timestamp 1704896540
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_43
timestamp 1704896540
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_13
timestamp 1704896540
transform 1 0 2300 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_36
timestamp 1704896540
transform 1 0 4416 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_34
timestamp 1704896540
transform 1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_40
timestamp 1704896540
transform 1 0 4784 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 1704896540
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1704896540
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_23
timestamp 1704896540
transform 1 0 3220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_36
timestamp 1704896540
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 1704896540
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1704896540
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1704896540
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1704896540
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_30
timestamp 1704896540
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_38
timestamp 1704896540
transform 1 0 4600 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_46
timestamp 1704896540
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1704896540
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1704896540
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1704896540
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704896540
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 in[0]
port 2 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 in[1]
port 3 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 in[2]
port 4 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 in[3]
port 5 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 in[4]
port 6 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 in[5]
port 7 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 in[6]
port 8 nsew signal input
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 in[7]
port 9 nsew signal input
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 480 0 0 0 out[0]
port 10 nsew signal output
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 480 0 0 0 out[1]
port 11 nsew signal output
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 480 0 0 0 out[2]
port 12 nsew signal output
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 480 0 0 0 out[3]
port 13 nsew signal output
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 480 0 0 0 out[4]
port 14 nsew signal output
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 480 0 0 0 out[5]
port 15 nsew signal output
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 480 0 0 0 out[6]
port 16 nsew signal output
flabel metal3 s 6100 824 6900 944 0 FreeSans 480 0 0 0 out[7]
port 17 nsew signal output
rlabel metal1 3450 8704 3450 8704 0 VGND
rlabel metal1 3450 9248 3450 9248 0 VPWR
rlabel metal1 4462 2890 4462 2890 0 _00_
rlabel metal1 3358 4590 3358 4590 0 _01_
rlabel metal2 4462 4114 4462 4114 0 _02_
rlabel metal1 4324 5542 4324 5542 0 _03_
rlabel metal1 3726 7174 3726 7174 0 _04_
rlabel metal1 4968 3162 4968 3162 0 _05_
rlabel metal1 3450 4114 3450 4114 0 _06_
rlabel via2 2070 4029 2070 4029 0 _07_
rlabel metal1 1656 4114 1656 4114 0 _08_
rlabel metal3 1050 10404 1050 10404 0 in[0]
rlabel metal3 751 9044 751 9044 0 in[1]
rlabel metal3 751 7684 751 7684 0 in[2]
rlabel metal3 751 6324 751 6324 0 in[3]
rlabel metal3 751 4964 751 4964 0 in[4]
rlabel metal3 751 3604 751 3604 0 in[5]
rlabel metal3 820 2244 820 2244 0 in[6]
rlabel metal3 1096 884 1096 884 0 in[7]
rlabel metal1 4324 5678 4324 5678 0 net1
rlabel metal1 4370 8874 4370 8874 0 net10
rlabel metal1 4094 4726 4094 4726 0 net11
rlabel metal1 3864 5134 3864 5134 0 net12
rlabel metal2 4370 4998 4370 4998 0 net13
rlabel metal2 5198 5134 5198 5134 0 net14
rlabel metal2 4646 2465 4646 2465 0 net15
rlabel metal2 5106 3162 5106 3162 0 net16
rlabel metal1 4508 5882 4508 5882 0 net2
rlabel metal2 3266 3774 3266 3774 0 net3
rlabel metal2 3174 5916 3174 5916 0 net4
rlabel metal2 4002 3468 4002 3468 0 net5
rlabel metal2 4094 3842 4094 3842 0 net6
rlabel metal1 2208 3978 2208 3978 0 net7
rlabel metal1 4692 4114 4692 4114 0 net8
rlabel metal1 4784 6426 4784 6426 0 net9
rlabel metal2 5014 9775 5014 9775 0 out[0]
rlabel via2 5382 9061 5382 9061 0 out[1]
rlabel via2 5382 7701 5382 7701 0 out[2]
rlabel metal2 5382 6477 5382 6477 0 out[3]
rlabel via2 5382 4981 5382 4981 0 out[4]
rlabel metal2 5382 3757 5382 3757 0 out[5]
rlabel via2 4830 2261 4830 2261 0 out[6]
rlabel metal2 5474 1615 5474 1615 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
